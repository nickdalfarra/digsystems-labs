library verilog;
use verilog.vl_types.all;
entity Bus32bit is
    port(
        i0out           : in     vl_logic;
        i1out           : in     vl_logic;
        i2out           : in     vl_logic;
        i3out           : in     vl_logic;
        i4out           : in     vl_logic;
        i5out           : in     vl_logic;
        i6out           : in     vl_logic;
        i7out           : in     vl_logic;
        i8out           : in     vl_logic;
        i9out           : in     vl_logic;
        i10out          : in     vl_logic;
        i11out          : in     vl_logic;
        i12out          : in     vl_logic;
        i13out          : in     vl_logic;
        i14out          : in     vl_logic;
        i15out          : in     vl_logic;
        i16out          : in     vl_logic;
        i17out          : in     vl_logic;
        i18out          : in     vl_logic;
        i19out          : in     vl_logic;
        i20out          : in     vl_logic;
        i21out          : in     vl_logic;
        i22out          : in     vl_logic;
        i23out          : in     vl_logic;
        i24out          : in     vl_logic;
        i25out          : in     vl_logic;
        i26out          : in     vl_logic;
        i27out          : in     vl_logic;
        i28out          : in     vl_logic;
        i29out          : in     vl_logic;
        i30out          : in     vl_logic;
        i31out          : in     vl_logic;
        i0              : in     vl_logic_vector(31 downto 0);
        i1              : in     vl_logic_vector(31 downto 0);
        i2              : in     vl_logic_vector(31 downto 0);
        i3              : in     vl_logic_vector(31 downto 0);
        i4              : in     vl_logic_vector(31 downto 0);
        i5              : in     vl_logic_vector(31 downto 0);
        i6              : in     vl_logic_vector(31 downto 0);
        i7              : in     vl_logic_vector(31 downto 0);
        i8              : in     vl_logic_vector(31 downto 0);
        i9              : in     vl_logic_vector(31 downto 0);
        i10             : in     vl_logic_vector(31 downto 0);
        i11             : in     vl_logic_vector(31 downto 0);
        i12             : in     vl_logic_vector(31 downto 0);
        i13             : in     vl_logic_vector(31 downto 0);
        i14             : in     vl_logic_vector(31 downto 0);
        i15             : in     vl_logic_vector(31 downto 0);
        i16             : in     vl_logic_vector(31 downto 0);
        i17             : in     vl_logic_vector(31 downto 0);
        i18             : in     vl_logic_vector(31 downto 0);
        i19             : in     vl_logic_vector(31 downto 0);
        i20             : in     vl_logic_vector(31 downto 0);
        i21             : in     vl_logic_vector(31 downto 0);
        i22             : in     vl_logic_vector(31 downto 0);
        i23             : in     vl_logic_vector(31 downto 0);
        i24             : in     vl_logic_vector(31 downto 0);
        i25             : in     vl_logic_vector(31 downto 0);
        i26             : in     vl_logic_vector(31 downto 0);
        i27             : in     vl_logic_vector(31 downto 0);
        i28             : in     vl_logic_vector(31 downto 0);
        i29             : in     vl_logic_vector(31 downto 0);
        i30             : in     vl_logic_vector(31 downto 0);
        i31             : in     vl_logic_vector(31 downto 0);
        busmux_out      : out    vl_logic_vector(31 downto 0)
    );
end Bus32bit;
