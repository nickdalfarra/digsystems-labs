library verilog;
use verilog.vl_types.all;
entity Datapath is
    port(
        Cout            : in     vl_logic;
        HIout           : in     vl_logic;
        LOout           : in     vl_logic;
        Zhighout        : in     vl_logic;
        Zlowout         : in     vl_logic;
        PCout           : in     vl_logic;
        MDRout          : in     vl_logic;
        BAout           : in     vl_logic;
        Inportout       : in     vl_logic;
        clear           : in     vl_logic;
        clk             : in     vl_logic;
        read            : in     vl_logic;
        write           : in     vl_logic;
        PCin            : in     vl_logic;
        IRin            : in     vl_logic;
        MARin           : in     vl_logic;
        Yin             : in     vl_logic;
        HIin            : in     vl_logic;
        LOin            : in     vl_logic;
        Zin             : in     vl_logic;
        MDRin           : in     vl_logic;
        Gra             : in     vl_logic;
        Grb             : in     vl_logic;
        Grc             : in     vl_logic;
        Rin             : in     vl_logic;
        Rout            : in     vl_logic;
        strobe          : in     vl_logic;
        OutPort         : in     vl_logic;
        \AND\           : in     vl_logic;
        \OR\            : in     vl_logic;
        ADD             : in     vl_logic;
        SUB             : in     vl_logic;
        MUL             : in     vl_logic;
        DIV             : in     vl_logic;
        SHR             : in     vl_logic;
        SHL             : in     vl_logic;
        \ROR\           : in     vl_logic;
        \ROL\           : in     vl_logic;
        NEG             : in     vl_logic;
        \NOT\           : in     vl_logic;
        IncPC           : in     vl_logic;
        CONin           : in     vl_logic;
        CON_FF          : out    vl_logic;
        InPortIn        : in     vl_logic_vector(31 downto 0);
        R0              : out    vl_logic_vector(31 downto 0);
        R1              : out    vl_logic_vector(31 downto 0);
        R2              : out    vl_logic_vector(31 downto 0);
        R3              : out    vl_logic_vector(31 downto 0);
        R4              : out    vl_logic_vector(31 downto 0);
        R5              : out    vl_logic_vector(31 downto 0);
        R6              : out    vl_logic_vector(31 downto 0);
        R7              : out    vl_logic_vector(31 downto 0);
        R8              : out    vl_logic_vector(31 downto 0);
        R9              : out    vl_logic_vector(31 downto 0);
        R10             : out    vl_logic_vector(31 downto 0);
        R11             : out    vl_logic_vector(31 downto 0);
        R12             : out    vl_logic_vector(31 downto 0);
        R13             : out    vl_logic_vector(31 downto 0);
        R14             : out    vl_logic_vector(31 downto 0);
        R15             : out    vl_logic_vector(31 downto 0);
        Hi              : out    vl_logic_vector(31 downto 0);
        Lo              : out    vl_logic_vector(31 downto 0);
        PC              : out    vl_logic_vector(31 downto 0);
        bus_mux_out     : out    vl_logic_vector(31 downto 0);
        IR              : out    vl_logic_vector(31 downto 0);
        MAR             : out    vl_logic_vector(31 downto 0);
        C_sign_ext      : out    vl_logic_vector(31 downto 0);
        InPortOutput    : out    vl_logic_vector(31 downto 0);
        OutPortOut      : out    vl_logic_vector(31 downto 0);
        Mdatain         : out    vl_logic_vector(31 downto 0);
        MDR             : out    vl_logic_vector(31 downto 0);
        Z               : out    vl_logic_vector(63 downto 0);
        ALUout          : out    vl_logic_vector(63 downto 0);
        Rins            : out    vl_logic_vector(15 downto 0);
        Routs           : out    vl_logic_vector(15 downto 0);
        ram_data        : inout  vl_logic_vector(31 downto 0);
        test1           : out    vl_logic;
        test2           : out    vl_logic;
        test3           : out    vl_logic;
        test4           : out    vl_logic
    );
end Datapath;
