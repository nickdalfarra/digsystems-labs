library verilog;
use verilog.vl_types.all;
entity Adder2bit_tb is
end Adder2bit_tb;
