library verilog;
use verilog.vl_types.all;
entity Divider32bit_tb is
end Divider32bit_tb;
