library verilog;
use verilog.vl_types.all;
entity MDR_tb is
end MDR_tb;
