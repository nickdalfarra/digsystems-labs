library verilog;
use verilog.vl_types.all;
entity conff_logic_tb is
end conff_logic_tb;
