library verilog;
use verilog.vl_types.all;
entity Bus32bit_tb is
end Bus32bit_tb;
