module Mux32bit32to1(input [4:0] select, input [31:0] i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, i22, i23, i24, i25, i26, i27, i28, i29, i30, i31, output [31:0] out);
	
	Mux8bit32to1 mux1 (select, i0[31:24], i1[31:24], i2[31:24], i3[31:24], i4[31:24], i5[31:24], i6[31:24], i7[31:24], i8[31:24], i9[31:24], i10[31:24], i11[31:24], i12[31:24], i13[31:24], i14[31:24], i15[31:24], i16[31:24], i17[31:24], i18[31:24], i19[31:24], i20[31:24], i21[31:24], i22[31:24], i23[31:24], i24[31:24], i25[31:24], i26[31:24], i27[31:24], i28[31:24], i29[31:24], i30[31:24], i31[31:24], out[31:24]);
	Mux8bit32to1 mux2 (select, i0[23:16], i1[23:16], i2[23:16], i3[23:16], i4[23:16], i5[23:16], i6[23:16], i7[23:16], i8[23:16], i9[23:16], i10[23:16], i11[23:16], i12[23:16], i13[23:16], i14[23:16], i15[23:16], i16[23:16], i17[23:16], i18[23:16], i19[23:16], i20[23:16], i21[23:16], i22[23:16], i23[23:16], i24[23:16], i25[23:16], i26[23:16], i27[23:16], i28[23:16], i29[23:16], i30[23:16], i31[23:16], out[23:16]);
	Mux8bit32to1 mux3 (select, i0[15:8], i1[15:8], i2[15:8], i3[15:8], i4[15:8], i5[15:8], i6[15:8], i7[15:8], i8[15:8], i9[15:8], i10[15:8], i11[15:8], i12[15:8], i13[15:8], i14[15:8], i15[15:8], i16[15:8], i17[15:8], i18[15:8], i19[15:8], i20[15:8], i21[15:8], i22[15:8], i23[15:8], i24[15:8], i25[15:8], i26[15:8], i27[15:8], i28[15:8], i29[15:8], i30[15:8], i31[15:8], out[15:8]);
	Mux8bit32to1 mux4 (select, i0[7:0], i1[7:0], i2[7:0], i3[7:0], i4[7:0], i5[7:0], i6[7:0], i7[7:0], i8[7:0], i9[7:0], i10[7:0], i11[7:0], i12[7:0], i13[7:0], i14[7:0], i15[7:0], i16[7:0], i17[7:0], i18[7:0], i19[7:0], i20[7:0], i21[7:0], i22[7:0], i23[7:0], i24[7:0], i25[7:0], i26[7:0], i27[7:0], i28[7:0], i29[7:0], i30[7:0], i31[7:0], out[7:0]);
	
endmodule
