library verilog;
use verilog.vl_types.all;
entity Encoder32to5 is
    port(
        i0              : in     vl_logic;
        i1              : in     vl_logic;
        i2              : in     vl_logic;
        i3              : in     vl_logic;
        i4              : in     vl_logic;
        i5              : in     vl_logic;
        i6              : in     vl_logic;
        i7              : in     vl_logic;
        i8              : in     vl_logic;
        i9              : in     vl_logic;
        i10             : in     vl_logic;
        i11             : in     vl_logic;
        i12             : in     vl_logic;
        i13             : in     vl_logic;
        i14             : in     vl_logic;
        i15             : in     vl_logic;
        i16             : in     vl_logic;
        i17             : in     vl_logic;
        i18             : in     vl_logic;
        i19             : in     vl_logic;
        i20             : in     vl_logic;
        i21             : in     vl_logic;
        i22             : in     vl_logic;
        i23             : in     vl_logic;
        i24             : in     vl_logic;
        i25             : in     vl_logic;
        i26             : in     vl_logic;
        i27             : in     vl_logic;
        i28             : in     vl_logic;
        i29             : in     vl_logic;
        i30             : in     vl_logic;
        i31             : in     vl_logic;
        \out\           : out    vl_logic_vector(4 downto 0)
    );
end Encoder32to5;
